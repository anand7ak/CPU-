
package test_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "half_adder_transaction.sv"
`include "half_adder_driver.sv"
`include "half_adder_monitor.sv"
`include "half_adder_scoreboard.sv"
`include "half_adder_agent.sv"
`include "half_adder_env.sv"
`include "test.sv"

endpackage
